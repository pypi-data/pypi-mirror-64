rc circuit

* pingspice:
* Object-oriented circuit construction and efficient asynchronous
* simulation with Ngspice and twisted.
*
* Copyright (C) 2017 by Edwin A. Suominen,
* http://edsuom.com/pingspice
*
* See edsuom.com for API documentation as well as information about
* Ed's background and other projects, software and otherwise.
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the
* License. You may obtain a copy of the License at
*
*   http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing,
* software distributed under the License is distributed on an "AS
* IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either
* express or implied. See the License for the specific language
* governing permissions and limitations under the License.

* Simple illustration of the RC time constant
* with big high-current components
* -------------------------------------------------------
* Deep-cycle battery
V1 1 0 dc 12 ac 1 PULSE(0, 12, 0, 1E-6)
* Wire series resistance
R1 1 2 0.1

* Big electrolytic capacitor to ground with 16 mOhm ESR
* and 20nH self-inductance
C1 2 3 47000u ic=0
R2 3 4 0.016
L2 4 0 20n

* A DC load that only turns on with enough voltage, and uses one extra
* amp for each extra volt it sees
R3 2 5 1
A1 0 5 turnon
.model turnon zener(v_breakdown=8.0, i_breakdown=1.0)

.CONTROL
set nomoremode
option reltol=0.01
option abstol=1e-09
option trtol=3.0
option gmin=1e-10
option itl4=20
option trytocompact
option vntol=1e-05
option itl1=200
option method=gear
option chgtol=1e-11
.ENDC

.END
