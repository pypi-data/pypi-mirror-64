.title Resistor Bridge
Vinput 1 0 10V
R1 1 2 2
R2 1 3 1
R3 2 0 1
R4 3 0 2
R5 3 2 2
** .op
* analysis 1
*.dc Vinput 10 20 1
*.save v(2) v(1)
* analysis 2
.sens v(1)
.end

