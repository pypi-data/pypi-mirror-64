OPAMP2.CIR - OPAMP MODEL (LEVEL 2)
* from http://www.ecircuitcenter.com/OpModels/OpampModels.htm
*
* SIGNAL SOURCE
VS	1	0	AC 1	PWL(0US 0V   0.01US 1V  100US 1V)
*
* POWER SUPPLIES
VCC	10	0	DC	+15V
VEE	11	0	DC	-15V
*
R1	0	2	1
*R2	2	3	1
XOP	1 2 3  10 11	OPAMP2
RL	3	0	100K
*
*
* OPAMP MACRO MODEL (INTERMEDIATE LEVEL)
*
*                IN+ IN- OUT  VCC  VEE
.SUBCKT OPAMP2   1   2   81   101   102  
Q1	5 1	7	NPN
Q2	6 2	8	NPN
RC1	101	5	95.49
RC2	101	6	95.49
RE1	7	4	43.79
RE2	8	4	43.79
I1	4	102	0.001
*
* OPEN-LOOP GAIN, FIRST POLE AND SLEW RATE
G1	100 10	6 5 0.0104719
RP1	10	100	9.549MEG
CP1	10	100	0.0016667UF
*
*OUTPUT STAGE
EOUT	80 100	10 100	1
RO	80	81	100
*
* INTERNAL REFERENCE
RREF1	101	103	100K
RREF2	103	102	100K
EREF	100 0	103 0 1
R100	100	0	1MEG
*
.model NPN  NPN(BF=50000)
*
.ENDS
*
* ANALYSIS
.TRAN 	0.1US  5US
.AC 	DEC 	5 0.1HZ 10MEGHZ
*
* VIEW RESULTS
.PRINT	TRAN 	V(3)
.PRINT	AC 	V(3)
.PROBE
.END
